module FSM (

);




endmodule 