`timescale 1 ps / 1 ps

module ir_controller_tb;

    // Testbench signals
    logic clk;
    logic rst_n;
    logic [31:0] ir_data;
    logic data_ready;
    logic drive, stop, increase_speed, decrease_speed, turn_left, turn_right;

    // Instantiate the ir_controller module
    ir_controller dut (
        .clk(clk),
        .rst_n(rst_n),
        .ir_data(ir_data),
        .data_ready(data_ready),
        .drive(drive),
        .stop(stop),
        .increase_speed(increase_speed),
        .decrease_speed(decrease_speed),
        .turn_left(turn_left),
        .turn_right(turn_right)
    );

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 10 ps clock period
    end

    // Test procedure
    initial begin
        // Reset the system
        rst_n = 0;
        #10 rst_n = 1;

        // Test the Power button (drive command)
        ir_data = 32'h00000012; // 0x12 is the key code for the power button
        data_ready = 1;
        #10 data_ready = 0;
        #10 $display("Drive: %b", drive); // Should print 1

        // Test the Mute button (stop command)
        ir_data = 32'h0000000C; // 0x0C is the key code for the mute button
        data_ready = 1;
        #10 data_ready = 0;
        #10 $display("Stop: %b", stop); // Should print 1

        // Test Volume Up (increase speed)
        ir_data = 32'h0000001B; // 0x1B is the key code for volume up
        data_ready = 1;
        #10 data_ready = 0;
        #10 $display("Increase Speed: %b", increase_speed); // Should print 1

        // Test Volume Down (decrease speed)
        ir_data = 32'h0000001F; // 0x1F is the key code for volume down
        data_ready = 1;
        #10 data_ready = 0;
        #10 $display("Decrease Speed: %b", decrease_speed); // Should print 1

        // Test Left Arrow (turn left)
        ir_data = 32'h00000014; // 0x14 is the key code for the left arrow
        data_ready = 1;
        #10 data_ready = 0;
        #10 $display("Turn Left: %b", turn_left); // Should print 1

        // Test Right Arrow (turn right)
        ir_data = 32'h00000018; // 0x18 is the key code for the right arrow
        data_ready = 1;
        #10 data_ready = 0;
        #10 $display("Turn Right: %b", turn_right); // Should print 1

        $stop; // End simulation
    end

endmodule

