module FSM (

);

endmodule 